boot02  hobgzhur.cre| Boots of Stealth             | hobgoblin from Zhurlong quest
                    |                              | 
brac07  hairto.cre  | Gauntlets of Dexterity       | Hairtooth, ogrillon near the gnoll stronghold
brac10  meilum.cre  | Gauntlets of Weapon Expertise| Meilum, the Sword Coast's most skilled swordsman
brac04  zal.cre     | Bracers of Archery           | Zal, the fastest dart thower
                    |                              | 
clck03  ulgoth.sto  | Cloak of Displacement        | store in Ulgoth's Beard
clck07  halbaz.dlg  | Nymph Cloak                  | Halbazzer Drin, Sorcerous Sundries
clck07  halbaz.cre  | Nymph Cloak                  | Halbazzer Drin, Sorcerous Sundries
clck15  highhedg.sto| Robe of the Good Archmagi    | High Hedge mage shop
clck16  highhedg.sto| Robe of the Neutral Archmagi | High Hedge mage shop
clck17  davaeo.cre  | Robe of the Evil Archmagi    | Davaeorn (BG1 mage who rules mines)
                    |                              | 
ring21  nimbul.cre  | Ring of Infravision          | Nimbul (asassin in Nashkel)
ring22  mulahe.cre  | Ring of Holiness             | Mulahey
