amul01  trcar04.sto                    | Necklace of Missiles           | merchant in Trademeet
amul16  ar0602.are                     | Metaspell Influence Amulet     | Jon's dungeon (container 11)
amul20  uddrow24.sto                   | Kaligun's Amulet of Magic Res. | Ust Natha store
amul21  aran02.cre                     | Amulet of Power                | Aran Linvail (side with Bodhi)
amul21  aran.dlg                       | Amulet of Power                | Aran Linvail (side with thieves)
amul24  ar0705.are                     | Necklace of Form Stability     | Merkath's lab (container 8)
regisamu c6regis.cre                   | Ruby Pendant                   | Regis (Drizzt's party)
regisamu c6regis2.cre                  | Ruby Pendant                   | Regis (Drizzt's party)
                                       |                                | 
belt02  mgkhol01.dlg                   | Golden Girdle                  | Sphere, Solamnic Knights, Khollynnus Paac
belt03  ar0603.are                     | Girdle of Bluntness            | Jon's dungeon lvl 2 (container 1)
belt04  kalah2.cre                     | Girdle of Piercing             | Kalah - circus
belt07  suadsaan.cre                   | Girdle of Stone Giant Strength | Suldanessellar Adsaan
belt09  gaal01.cre                     | Girdle of Fortitude            | Cult of Eyeless, Gaal
                                       |                                | 
boot03  tokcre01.dlg                   | Boots of the North             | Token machine in Spellhold
boot05  tokcre01.dlg                   | Boots of Grounding             | Token machine in Spellhold
boot04  reti.cre                       | Boots of Avoidance             | Reti (Buried alive quest)
boot11  ar2300.are                     | Boots of Etherealness          | Sahuagin city (chest 6)
boot12  amsmug02.sto                   | Gargoyle Boots                 | Carras, Amekthran smuggler
                                       |                                | 
brac03  lyros.cre                      | Bracers of Defense AC 6        | Xzar (Harpers quest)
brac06  obshal01.cre                   | Gauntlets of Ogre Power        | Lavok's sphere, Entu
brac09  pthral05.cre                   | Gauntlets of Weapon Skill      | Planar Prison, Female Thrall (Haerdalis quest)
brac14  udsvir05.dlg                   | Bracers of Defense AC 4        | Underdark, svirf innkeeper (reward for rescuing his son)
brac15  ribald.sto                     | Bracers of Defense AC 3        | Ribald
brac16  udprince.cre                   | Bracers of Blinding Strike     | Underdark, Kuo-Toa Prince
brac18  trthf01.cre                    | Gloves of Missile Snaring      | Itona the Shadow Thief in Trademeet
brac19  sahkng01.dlg                   | Gauntlets of Crushing          | Sahuagin city, King Ixilthetocal
brac21  gorwom03.cre                   | Gauntlets of Extraordinary Spec| Watcher's Keep last level, Y'tossi
brac26  bazdra02.cre                   | Tzu-Zan's Bracers              | Draconis
                                       |                                | 
clck06  sevpat02.cre                   | Cloak of Non-Detection         | Sorcerous Amon (Seven Vales party)
clck24  ar1511.are                     | Cloak of Reflection            | Spellhold (container 1)
clck27  sewrak01.cre                   | Cloak of the Sewers            | Rakshasa in sewers
clck04  shabod01.cre                   | Cloak of the Wolf              | Wallag's body (no idea who is this)
                                       |                                | 
ring02  firrak01.cre                   | Ring of Fire Resistance        | rakshasa in Firkraag's lair
ring04  ar2210.are                     | Ring of Clumsiness             | Ust Natha, lich tower
ring05  grvlch01.cre                   | Ring of Invisibility           | lich at City Gates
ring08  ar0411.bcs                     | Ring of Wizardry, BG2 version  | mage stronghold (if all apprentices die)
ring08  mgappr02.dlg                   | Ring of Wizardry, BG2 version  | mage stronghold (if Morul lives)
ring09  ppbook.bcs                     | Ring of Free Action            | book on the stand in spellhold
ring20  ribald.sto                     | Ring of Energy                 | Ribald
ring23  ar2100.are                     | Ring of Folly                  | Underdark svirf village (container 6)
ring30  kalah2.cre                     | Ring of Human Influence        | Kalah - circus
ring31  ppstat01.dlg                   | Ring of Regeneration           | statue in Spellhold
ring34  udardul.cre                    | Ring of Spell Turning          | Underdark, matron mother Ardulace
ring35  arnman09.cre                   | Ring of Lock Picks             | Shadow thieves, we're with Aran
ring35  arnwar07.cre                   | Ring of Lock Picks             | Shadow thieves, we're with Bodhi
ring36  ar0413.are                     | Ring of Danger Sense           | Planar Sphere container 1
ring39  hldemi.cre                     | Ring of Gaxx                   | Kangaxx
ring42  bazdra03.cre                   | Ring of Improved Invisibility  | Fll'Yissetat Abazigal's dragon-guard
// ring43 is RoP+3 from deck - skipping|                                | 
                                       |                                | 
helm04  hlmafer.cre                    | Helm Of Defence                | Maferan (Guarded compound)
dagg03  c6arkan.cre                    | Dagger +2: 'Heart of the Golem'| Arcanis Gath in Bodhi's lair (1 and 2 stage, possibly)
dagg03  c6arkan3.cre                   | Dagger +2: 'Heart of the Golem'| Arcanis Gath in Bodhi's lair (1 and 2 stage, possibly)
shld19  chak.cre                       | Large Shield +2                | Chak (Firkraag's dungeon, Samia's party)
sw1h10  renal.cre                      | Short Sword of Backstabbing +3 | Renal Bloodscalp
sw1h10  renal.dlg                      | Short Sword of Backstabbing +3 | Renal Bloodscalp
halb03  jarevia.cre                    | Suryris's Blade                | Reviane - Jaheira's quest
sw1h03  lehtin.dlg                     | Kondar +1, +3 vs Shapeshifters | Lehtinan (Copper coronet)
sw1h03  hendak.dlg                     | Kondar +1, +3 vs Shapeshifters | Hendak (Copper coronet)
sw1h06  ribald.cre                     | Long Sword +2: 'Varscona'      | Ribald - both EE and fixpack ensure it's unique
wa2robe wmart2.sto                     | Robe of Vecna                  | Deidre
