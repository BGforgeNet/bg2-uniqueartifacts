amul14  nadine.cre                       | Necklace of Missiles           | Nadine - steal
amul14  nadin.dlg                        | Necklace of Missiles           | Nadine - quest reward
amul16  ramazi.cre                       | Metaspell Influence Amul.      | Ramazith
                                         |                                | 
belt02  kirian.cre                       | Golden Girdle                  | Kirian - band in Mutamin's garden
belt03  krumm.cre                        | Girdle of Bluntness            | the guy who cuts nymph's tree
belt04  ogreunsh.cre                     | Girdle of Piercing             | fetishist ogre
                                         |                                | 
boot03  jared.cre                        | Boots of the North             | Jared the scared merchant (a bear and a bridge) - steal
boot03  jared.dlg                        | Boots of the North             | Jared the scared merchant (a bear and a bridge) - talk
boot04  nimbul.cre                       | Boots of Avoidance             | Nimbul, assassin in Nashkel
boot05  mulahe.cre                       | Boots of Grounding             | Mulahey
                                         |                                | 
brac03  davaeo.cre                       | Bracers of Defense AC 6        | Davaeorn - Cloakwood mines boss
brac06  desret.cre                       | Gauntlets of Ogre Power        | Desreta, assasin in tavern-ship
brac08  bassil.cre                       | Gauntlets of Fumbling          | Bassilus - BG1 only, not present in BG2
brac09  %BaldursGateDocks%.are           | Gauntlets of Weapon Skill      | BG docks, chest near Umberlee temple (Noralee's quest)
                                         |                                | 
clck04  %Lighthouse_BlackAlaricsCave%.are| Cloak of the Wolf              | Black Alarick's Cave
clck05  quenas.cre                       | Cloak of Balduran              | Quenash - steal
clck05  quenas.dlg                       | Cloak of Balduran              | Quenash - talk
clck06  taslgurk.cre                     | Cloak of Non-Detection         | Gurke's tasloi, Cloakwood 1
clck08  algern.cre                       | Algernon's Cloak               | Algernon, Beregost
                                         |                                | 
ring02  %Candlekeep_Catacombs_L1%.are    | Ring of Fire Resistance        | Candlekeep catacombs level 1
ring04  niemai.cre                       | Ring of Clumsiness             | Niemain, Sorcerous Sundries 2nd floor
ring05  ulgoth.sto                       | Ring of Invisibility           | store in Ulgoth's Beard
ring09  alai.cre                         | Ring of Free Action            | Alai, party at the top of the Iron Throne
ring20  denak.cre                        | Ring of Energy                 | Thaivian red wizard
ring23  %ShipwrecksCoast%.are            | Ring of Folly                  | shipwreck on the coast (container 1)
misc72  highhedg.sto                     | Claw of Kazgaroth              | when importing from BG1, may be found in import03.2da
                                         |                                | 
dagg03  hentol.cre                       | Dagger +2: 'Heart of the Golem'| Hentold in Valley of Tombs (give dagger to revenant)
dagg03  hentol.dlg                       | Dagger +2: 'Heart of the Golem'| Hentold in Valley of Tombs (give dagger to revenant)
halb03  zhalim.cre                       | Suryris's Blade                | party on the last level of Iron throne
helm04  droth.cre                        | Helmet of Defence                | Droth the ogre-mage who mates with a sirene
leat03  maneir.cre                       | Protector of the second        | Maneira, bounty hunters party
sw1h06  greywo.cre                       | Long Sword +2: 'Varscona'      | Greywolf (bounty hunter coming for Prism)
sw1h03  aldeth.cre                       | Kondar +1, +3 vs Shapeshifters | Aldeth Sashenstar (Cloakwood or BG) - should be droppable but not stealable, handled in custom.tpa
sw1h03  aldeth.dlg                       | Kondar +1, +3 vs Shapeshifters | Aldeth Sashenstar (Cloakwood or BG) - quest reward
sw1h10  slythe.cre                       | Short Sword of Backstabbing    | Slythe - last asassination attempt in underground tavern
