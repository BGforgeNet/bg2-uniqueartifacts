amul22  trrak01.cre | Periart of Proof against Poison  | Adratha/Ithafeer
amul23  scsain.dlg  | Periart of Life Protection       | Cleric of Lathander quest reward (stronghold illitium)
amul26  senken01.cre| Amulet of Cheetah Speed          | drow in Sendai enclave
amul28  elemimix.cre| Amulet of the Master Harper      | Imix - Yaga-Shura Castle
wa2amu  wmart2.sto  | Sensate Amulet                   | Deidre
                    |                                  | 
belt06  ribald.sto  | Girdle of Hill Giant Strength    | Ribald
belt08  uddeath2.cre| Girdle of Frost Giant Strength   | Underdark, Demon Knight
belt10  trmer02.sto | Belt of Inertial Barrier         | Merchant in Trademeet
belt11  ar5201.are  | Girdle of Fire Giant Strength    | 1st part Yaga-Shura's hold container 3
                    |                                  | 
boot02  ar0303.are  | Boots of Stealth                 | Maevar's Guild (container 5)
                    |                                  | 
brac04  ar1904.are  | Bracers of Archery               | troll mound near druid grove, container 2
brac07  ar0206.are  | Gauntlets of Dexterity           | Undead town, cont 1 (eyeless quest)
brac10  ar0808.are  | Gauntlets of Weapon Expertise    | 6th chapter, container 6
brac13  elelev01.dlg| Bracers of Defense AC 5          | machine in Spellhold
brac20  kayl2.dlg   | Gloves of Healing                | Sir Ryan Trawl quest reward
brac22  ar3001.are  | Paladin's Bracers                | Watcher's Keep 1st level, chest1
                    |                                  | 
clck03  trmer02.sto | Cloak of Displacement            | Merchant in Trademeet
clck07  gorch.sto   | Nymph Cloak                      | merchant Gorch in Maevar's guild
clck15  25spell.sto | Robe of the Good Archmagi        | Lazarus store in Saradush - ToB
clck15  trmer04.sto | Robe of the Good Archmagi        | Merchant in Trademeet
clck16  ribald2.sto | Robe of the Neutral Archmagi     | Ribald's enhanced shop
clck17  uddrow23.sto| Robe of the Evil Archmagi        | Ust Natha's shop
clck25  uhrang01.cre| Cloak of the Stars               | Merella
clck26  sahramb3.cre| Cloak of Mirroring               | sahuagin priestess
clck30  hellfear.dlg| Cloak of Bravery                 | hell trials, Fear
                    |                                  | 
ring03  govwau01.sto| Ring of Animal Friendship        | Waukeen temple in government district
ring22  alphonse.bcs| Ring of Holiness                 | Reward for illithium quest
ring26  ar0329.are  | Ring of Djinni Summoning         | Aran's guild (cont8), only available when siding with Bodhi
ring27  uddwarf.cre | Ring of Fire Control             | Mad dwarf in illithid lair in Underdark
ring28  ribald.sto  | Ring of Air Control              | Ribald
ring29  ar1302.are  | Ring of Earth Control            | De'Arnise Hold 1st floor container1
ring40  lavok01.cre | Ring of Acuity                   | Lavok
ring40  lavok02.cre | Ring of Acuity                   | Lavok
ring46  amlich01.cre| Ring of Anti-Venom               | Vongoethe (lich in ToB)
wa2ring  wmart2.sto | Mercykiller Ring                 | Deidre
                    |                                  | 
shld30  hlmafer.cre | Large Shield +2 - Calimport mercs| Maferan (Guarded compound)
sw1h53  bernard2.sto| Sword of Flame +1                | Bernard, after freeing slaves
xbow06  bernard2.sto| Light Crossbow of Speed          | Bernard, after freeing slaves
