wand02  ar1803.are  | Wand of Fear             | Cloakwood Mines, locked chest in Davaeorn's lair, 15 charges
wand02  beyn.cre    | Wand of Fear             | Beyn, fighter/mage on Ice Island, 13 charges
wand02  bpxith01.sto| Wand of Fear             | Xithiss, mind flayer merchant in Black Pits
wand02  bpxith02.sto| Wand of Fear             | Xithiss, mind flayer merchant in Black Pits
wand02  bpxith03.sto| Wand of Fear             | Xithiss, mind flayer merchant in Black Pits
wand02  highhedg.sto| Wand of Fear             | Thalantyr, mage shop in High Hedge, 20 charges
                    |                          | 
wand03  ar0603.are  | Wand of Magic Missiles   | Seven Suns, basement, 30 charges
wand03  ar1501.are  | Wand of Magic Missiles   | Balduran's ship, ground floor, 5 charges
wand03  bpxith01.sto| Wand of Magic Missiles   | Xithiss, mind flayer merchant in Black Pits
wand03  bpxith02.sto| Wand of Magic Missiles   | Xithiss, mind flayer merchant in Black Pits
wand03  bpxith03.sto| Wand of Magic Missiles   | Xithiss, mind flayer merchant in Black Pits
wand03  tranzi.cre  | Wand of Magic Missiles   | Tranzig, 2nd floor in Feldepost Inn, 31 charges
                    |                          | 
wand04  ar3601.are  | Wand of Paralyzation     | Black Alaric's cave, 13 charges
wand04  bpxith02.sto| Wand of Paralyzation     | Xithiss, mind flayer merchant in Black Pits
wand04  bpxith03.sto| Wand of Paralyzation     | Xithiss, mind flayer merchant in Black Pits
wand04  cuchol.cre  | Wand of Paralyzation     | Cuchol, fighter/mage on Ice Island, 11 charges
wand04  resar.cre   | Wand of Paralyzation     | Resar, Halruaan mage in Thieves' Guild, 12 charges
                    |                          | 
wand05  ar0514.are  | Wand of Fire             | Durlag's Tower, 5th subterranean level, 12 charges
wand05  ar2615.are  | Wand of Fire             | Candlekeep Catacombs, 1st level, 16 charges
wand05  ar3901.are  | Wand of Fire             | Ulcaster School, dungeon, 8 charges
wand05  bpxith01.sto| Wand of Fire             | Xithiss, mind flayer merchant in Black Pits
wand05  bpxith02.sto| Wand of Fire             | Xithiss, mind flayer merchant in Black Pits
wand05  bpxith03.sto| Wand of Fire             | Xithiss, mind flayer merchant in Black Pits
                    |                          | 
wand06  ar2101.are  | Wand of Frost            | Cloakwood, Spider Nest, 12 charges
wand06  ar5400.are  | Wand of Frost            | Nashkel Mines, tree, 10 charges
wand06  bpaluena.cre| Wand of Frost            | Thespia, ? in Black Pits
wand06  bpxith01.sto| Wand of Frost            | Xithiss, mind flayer merchant in Black Pits
wand06  bpxith02.sto| Wand of Frost            | Xithiss, mind flayer merchant in Black Pits
wand06  bpxith03.sto| Wand of Frost            | Xithiss, mind flayer merchant in Black Pits
wand06  centeo.cre  | Wand of Frost            | Centeol, Spider Nest in Cloakwood, undroppable
wand06  ulgoth.sto  | Wand of Frost            | Ulgoth's Beard, store, 29 charges
                    |                          | 
wand07  alai.cre    | Wand of Lightning        | Alai, party at the top of the Iron Throne, 10 charges
wand07  ar0504.are  | Wand of Lightning        | Durlag's Tower, third floor, 16 charges
wand07  ar3321.are  | Wand of Lightning        | Beregost, 2nd floor in Travenhurst Manor, 6 charges
wand07  bpxith01.sto| Wand of Lightning        | Xithiss, mind flayer merchant in Black Pits
wand07  bpxith02.sto| Wand of Lightning        | Xithiss, mind flayer merchant in Black Pits
wand07  bpxith03.sto| Wand of Lightning        | Xithiss, mind flayer merchant in Black Pits
                    |                          | 
wand08  cult2.cre   | Wand of Sleep            | Cult Wizard, Ulgoth's Beard, 4 charges
wand08  highhedg.sto| Wand of Sleep            | Thalantyr, mage shop in High Hedge, 20 charges
wand08  sto0703.sto | Wand of Sleep            | Halbazzer Drin, mage shop in Sorcerous Sundries, 20 charges
                    |                          | 
wand10  ar0511.are  | Wand of Monster Summoning| Durlag's Tower, second subterranean level, 5 charges
wand10  ar5001.are  | Wand of Monster Summoning| Valley of the Tombs, tomb, 8 charges
wand10  bpxith02.sto| Wand of Monster Summoning| Xithiss, mind flayer merchant in Black Pits
wand10  bpxith03.sto| Wand of Monster Summoning| Xithiss, mind flayer merchant in Black Pits
wand10  sto0703.sto | Wand of Monster Summoning| Halbazzer Drin, mage shop in Sorcerous Sundries, 20 charges
                    |                          | 
wand11  aasim.cre   | Wand of the Heavens      | Aasim, party at the top of the Iron Throne, 11 charges
wand11  bpxith03.sto| Wand of the Heavens      | Xithiss, mind flayer merchant in Black Pits
wand11  sto0703.sto | Wand of the Heavens      | Halbazzer Drin, mage shop in Sorcerous Sundries, 20 charges
wand11  ulgoth.sto  | Wand of the Heavens      | Ulgoth's Beard, store, 25 charges
